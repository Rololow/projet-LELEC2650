* TSMC 65nm Cascode Miller OTA Simulation - PSRR (Power Supply Rejection Ratio)
* December 2024
*-----------------------------------------------

************************************
*	Library & Technology settings
************************************

* Library containing the transistor model from the foundry
.LIB key=K1 '/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo' tt_lib

************************************
*	Include circuit definition
************************************

.include ./CascodeMillerOTA.cir

*******************************
*	Supply
*******************************

*** Supply voltage with AC for PSRR measurement
VVDD VDD GND DC vdd_val AC 1

*******************************
*	Stimuli - PSRR+ (positive supply)
*******************************

*** PSRR Measurement Setup
* Short inputs to ground (or DC bias)
* Apply AC signal on VDD
* Measure output response

.param V_IN_DC = 0.5

* Input bias (no AC, both inputs at same DC)
VVINp INp GND DC V_IN_DC
VVINm INm GND DC V_IN_DC

**********************************
*	Simulations
**********************************

.OP

*** AC analysis for PSRR
.param fmin = 1
.param fmax = 1Giga
.AC dec 100 fmin fmax

**********************************
*	Measurements
**********************************

*** Plot signals
.plot AC VDB(OUT) VP(OUT)

*** Supply to output gain (for PSRR calculation)
* PSRR = Adm / (Vout/Vdd) = Adm_dB - (Vout/Vdd)_dB

* Output response to supply variation
.extract AC label=Avdd_dB_1Hz 'yval(VDB(OUT),1)'
.extract AC label=Avdd_dB_1kHz 'yval(VDB(OUT),1e3)'
.extract AC label=Avdd_dB_1MHz 'yval(VDB(OUT),1e6)'
.extract AC label=Avdd_dB_max 'max(VDB(OUT))'

*** PSRR = Adm / Avdd = Adm_dB - Avdd_dB
* Using Adm from TB_AC (approximately 71.8 dB for this design)
.param Adm_dB = 71.8
.extract AC label=PSRR_1Hz 'Adm_dB - yval(VDB(OUT),1)'
.extract AC label=PSRR_1kHz 'Adm_dB - yval(VDB(OUT),1e3)'
.extract AC label=PSRR_1MHz 'Adm_dB - yval(VDB(OUT),1e6)'

*** DC operating point
.extract DC label=VOUT_DC V(OUT)
.extract DC label=Power '-V(VDD)*I(VVDD)'

.end
