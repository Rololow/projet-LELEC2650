* TSMC 65nm Miller OTA Simulation
* Sylvain Favresse & Grégoire Brandsteert
* November 2025
*-----------------------------------------------

*******************************
*	Options
*******************************

* Temperature
.temp 25

* To tune the accuracy of the simulation (related to the numerical methods, beyond the scope of this course; check the manual)
.option EPS = 1e-6

*******************************
* M1/M2: W = 1.77 um; L = 2.00 um
* M3/M4: W = 1.77 um; L = 2.00 um
* M5/M6: W = 0.48 um; L = 2.00 um
* M7/M8: W = 0.95 um; L = 2.00 um
* M9:    W = 17.70 um; L = 2.00 um
* M10:   W = 4.75 um; L = 2.00 um
* M11:   W = 3.54 um; L = 2.00 um
* M12:   W = 3.54 um; L = 2.00 um
* M13:   W = 0.95 um; L = 2.00 um
* M14:   W = 0.48 um; L = 2.00 um
* M15:   W = 0.48 um; L = 2.00 um
* IBIAS: 1.35 uA
* VIN MAX:   0.62 V
* VIN MIN:   -0.10 V
* VDSAT1:   0.15 V
* VIN:   0.26 V
* VOUT:  0.61 V
* Cf:    2.58 pF
*******************************

*** Supply voltage
.param vdd_val = 1.2

*** Load capacitance
.param Cl_val = 10p

*** Transistor dimensions - imported from sizing.cir
.include ./sizing.cir

*** AC simulation parameters

.param V0 = 5m
.param fmin = 1
.param fmax = 1e9
.param ac_dec = 20

*******************************
*	Device under test
*******************************

***** Miller OTA

* Reminder
* xMN D G S B


* netlist : 
* M14 VBIAS2 VBIAS2 0 0 NMOS
* M13 VBIAS3 VBIAS2 0 0 NMOS
* M15 VBIAS1 VBIAS1 VBIAS2 VBIAS2 NMOS
* M7 N007 VBIAS2 0 0 NMOS
* M8 N006 VBIAS2 0 0 NMOS
* M6 N001 VBIAS1 N007 N007 NMOS
* M5 N002 VBIAS1 N006 N006 NMOS
* M10 N003 VBIAS2 0 0 NMOS
* C1 N003 N002 Cm
* C2 N003 0 CL
* M4 N001 N001 VDD VDD PMOS
* M3 N002 N001 VDD VDD PMOS
* M9 N003 N002 VDD VDD PMOS
* M2 N006 VIN+ N005 N005 PMOS
* M1 N007 VIN- N005 N005 PMOS
* M11 N005 VBIAS3 VDD VDD PMOS
* M12 VBIAS3 VBIAS3 VDD VDD PMOS
* I1 VDD VBIAS1 I

xM1 N007 INm N005 N005 pch_lvt_mac W=W1 L=L1
xM2 N006 INp N005 N005 pch_lvt_mac W=W2 L=L2

xM3 N002 N001 VDD VDD pch_lvt_mac W=W3 L=L3
xM4 N001 N001 VDD VDD pch_lvt_mac W=W4 L=L4
xM5 N002 VBIAS1 N006 N006 nch_lvt_mac W=W5 L=L5
xM6 N001 VBIAS1 N007 N007 nch_lvt_mac W=W6 L=L6

xM7 N007 VBIAS2 GND GND nch_lvt_mac W=W7 L=L7
xM8 N006 VBIAS2 GND GND nch_lvt_mac W=W8 L=L8

xM9 OUT N002 VDD VDD pch_lvt_mac W=W9 L=L9
xM10 OUT VBIAS2 GND GND nch_lvt_mac W=W10 L=L10

xM11 N005 VBIAS3 VDD VDD pch_lvt_mac W=W11 L=L11
xM12 VBIAS3 VBIAS3 VDD VDD pch_lvt_mac W=W12 L=L12

xM13 VBIAS3 VBIAS2 GND GND nch_lvt_mac W=W13 L=L13
xM14  VBIAS2 VBIAS2 GND GND nch_lvt_mac W=W14 L=L14
xM15 VBIAS1 VBIAS1 VBIAS2 VBIAS2 nch_lvt_mac W=W15 L=L15
Cf OUT N002 Cf_val

* Load capacitance
Cload OUT GND Cl_val
	
**********************************
*	Supply and stimuli
**********************************

*** Ideal current source	
IIbias VDD VBIAS1 DC IBIAS

*** Ground
* absolute voltage reference
.connect GND 0

*** Supply voltage - DEFINED IN TESTBENCH
* VVDD VDD GND DC vdd_val