* TSMC 65nm Cascode Miller OTA Simulation - PVT Corners
* Based on TB_PVT.cir from TP6
* December 2024
*-----------------------------------------------

************************************
*	Library & Technology settings
************************************

* Library containing the transistor model from the foundry
.LIB key=K1 '/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo' tt_lib

************************************
*	Include circuit definition
************************************

.include ./CascodeMillerOTA.cir

*******************************
*	Supply
*******************************

*** Supply voltage
VVDD VDD GND DC vdd_val

*******************************
*	Stimuli
*******************************

*** Input Voltages Sources - Pseudo closed-loop operation
VSTB INm OUT
VVINp INP 0 DC VIN
.LSTB VSTB
*** See TP5 for more details


*******************************
*	PVT variations
*******************************

*** Temperature
.param temp_cold = -40
.param temp_hot = 85

*** Supply voltage (VDD0 = 1.2V from CascodeMillerOTA.cir)
.param VDD0 = 1.2
.param vdd_low = 0.9 * VDD0
.param vdd_high = 1.1 * VDD0


**********************************
*	Measurements
**********************************

.extract DC label=VINp V(INp)
.extract DC label=VINm V(INm)
.extract DC label=VOUT V(OUT)

*** Input pair M1/M2
.extract DC label=VGS1 VGS(xM1.MAIN)
.extract DC label=VDS1 VDS(xM1.MAIN)

*** Cascode transistors M5/M6
.extract DC label=VDS5 VDS(xM5.MAIN)
.extract DC label=VDS6 VDS(xM6.MAIN)

*** Output stage
.extract DC label=VSD9 -VDS(xM9.MAIN)
.extract DC label=VDS10 VDS(xM10.MAIN)

*** Currents
.extract DC label=ID1 I(xM1.MAIN.D)
.extract DC label=gm_over_ID1 'gm(xM1.MAIN)/ID1'
.extract DC label=Power '-V(VDD)*I(VVDD)'

* Region of operation
.extract DC label=M1 opmode(xM1.MAIN)
.extract DC label=M2 opmode(xM2.MAIN)
.extract DC label=M3 opmode(xM3.MAIN)
.extract DC label=M4 opmode(xM4.MAIN)
.extract DC label=M5 opmode(xM5.MAIN)
.extract DC label=M6 opmode(xM6.MAIN)
.extract DC label=M7 opmode(xM7.MAIN)
.extract DC label=M8 opmode(xM8.MAIN)
.extract DC label=M9 opmode(xM9.MAIN)
.extract DC label=M10 opmode(xM10.MAIN)
.extract DC label=M11 opmode(xM11.MAIN)
.extract DC label=M12 opmode(xM12.MAIN)
.extract DC label=M13 opmode(xM13.MAIN)
.extract DC label=M14 opmode(xM14.MAIN)
.extract DC label=M15 opmode(xM15.MAIN)

.extract DC label=gdeq 'GDS(xM9.MAIN)+GDS(xM10.MAIN)'

.extract DC label=gm1 gm(xM1.MAIN)
.extract DC label=gm9 gm(xM9.MAIN)
.extract DC label=Vth1 Vth(xM1.MAIN)

*** Gain

.plot AC LSTB_DB LSTB_P

* magnitude in dB
.extract AC label=Av0dB 'max(LSTB_DB)'
* absolute magnitude
.extract AC label=Av0 '10^(Av0dB/20)'

*** Transition Frequency
* Real value from AC simulation
.extract AC label=fT 'xthres(LSTB_DB,0)'

.extract AC label=Phase_Margin '180 - yval(LSTB_P,1) + xycond(LSTB_P,LSTB_DB<0)'

**********************************
*	Simulations
**********************************

.OP

.param fmin = 1
.param fmax = 1Giga
.AC dec 100 fmin fmax

*** Print PVT results to file (one line per corner)
.printfile AC meas(Av0dB) meas(Av0) meas(fT) meas(Phase_Margin) meas(Power) file=PVT_results.txt format=data


***** PVT corners - DC and AC *****


.alter FF_LOW_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ff_lib
.param vdd_val = vdd_low
.param temperature_val = temp_cold

.alter FF_LOW_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ff_lib
.param vdd_val = vdd_low
.param temperature_val = temp_hot

.alter FF_HIGH_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ff_lib
.param vdd_val = vdd_high
.param temperature_val = temp_cold

.alter FF_HIGH_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ff_lib
.param vdd_val = vdd_high
.param temperature_val = temp_hot

.alter SS_LOW_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ss_lib
.param vdd_val = vdd_low
.param temperature_val = temp_cold

.alter SS_LOW_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ss_lib
.param vdd_val = vdd_low
.param temperature_val = temp_hot

.alter SS_HIGH_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ss_lib
.param vdd_val = vdd_high
.param temperature_val = temp_cold

.alter SS_HIGH_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" ss_lib
.param vdd_val = vdd_high
.param temperature_val = temp_hot

.alter SF_LOW_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" sf_lib
.param vdd_val = vdd_low
.param temperature_val = temp_cold

.alter SF_LOW_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" sf_lib
.param vdd_val = vdd_low
.param temperature_val = temp_hot

.alter SF_HIGH_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" sf_lib
.param vdd_val = vdd_high
.param temperature_val = temp_cold

.alter SF_HIGH_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" sf_lib
.param vdd_val = vdd_high
.param temperature_val = temp_hot

.alter FS_LOW_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" fs_lib
.param vdd_val = vdd_low
.param temperature_val = temp_cold

.alter FS_LOW_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" fs_lib
.param vdd_val = vdd_low
.param temperature_val = temp_hot

.alter FS_HIGH_COLD
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" fs_lib
.param vdd_val = vdd_high
.param temperature_val = temp_cold

.alter FS_HIGH_HOT
.LIB key=K1 "/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo" fs_lib
.param vdd_val = vdd_high
.param temperature_val = temp_hot

.end
