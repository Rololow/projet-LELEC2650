* TSMC 65nm Cascode Miller OTA Simulation - CMRR (Common Mode Rejection Ratio)
* December 2024
*-----------------------------------------------

************************************
*	Library & Technology settings
************************************

* Library containing the transistor model from the foundry
.LIB key=K1 '/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo' tt_lib

************************************
*	Include circuit definition
************************************

.include ./CascodeMillerOTA.cir

*******************************
*	Supply
*******************************

*** Supply voltage
VVDD VDD GND DC vdd_val

*******************************
*	Stimuli
*******************************

*** CMRR Measurement Setup
* Apply same AC signal to both inputs (common mode)
* Measure output response

.param V_CM_DC = VIN
.param V_AC = 1m

* Common mode input: same signal on both inputs
VVINp INp GND DC V_CM_DC AC V_AC
VVINm INm GND DC V_CM_DC AC V_AC

**********************************
*	Simulations
**********************************

.OP

*** AC analysis for common mode gain
* Use the global AC parameters from the device include so all TBs share the same grid
.AC dec ac_dec fmin fmax

**********************************
*	Measurements
**********************************

*** Plot signals
.plot AC VDB(OUT) VP(OUT)

*** Common mode gain (Acm)
.extract AC label=Acm_dB_1Hz 'yval(VDB(OUT),1)'
.extract AC label=Acm_dB_1kHz 'yval(VDB(OUT),1e3)'
.extract AC label=Acm_dB_1MHz 'yval(VDB(OUT),1e6)'
.extract AC label=Acm_dB_max 'max(VDB(OUT))'

*** Note: CMRR will be computed in python by subtracting cm_gain (this file)
*** from the differential gain exported by `TB_AC.cir` (diff_gain.txt).

*** DC operating point
.extract DC label=VOUT_DC V(OUT)
.extract DC label=Power '-V(VDD)*I(VVDD)'

* ------------------------------------------------------------------
* Example export (ASCII) for common-mode gain (frequency, Av_cm_dB)
* Uncomment to write `cm_gain.txt` which `plot_results.py` can read.
* Syntax may vary with Eldo versions; adjust if needed.
*
.printfile AC VDB(OUT) file=cm_gain.txt format=data
*
* To create the differential gain file, run `TB_AC.cir` (differential stimulus)
* and enable the diff export in that TB (see diff_gain.txt example there).
* ------------------------------------------------------------------

.end
