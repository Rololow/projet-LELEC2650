* TSMC 65nm Miller OTA Simulation
* Sylvain Favresse & Grégoire Brandsteert
* November 2025
*-----------------------------------------------

************************************
*	Library & Technology settings
************************************

* Library containing the transistor model from the foundry
.lib '/dir/TECHNOLOGY/cds2024/TSMC-N65/CMOS/LP/pdk/models/eldo/toplevel.eldo' tt_lib

*******************************
*	Options
*******************************

* Temperature
.temp 25

* To tune the accuracy of the simulation (related to the numerical methods, beyond the scope of this course; check the manual)
.option EPS = 1e-6

*******************************
* M1/M2: W = 3.18 um; L = 2.00 um
* M3/M4: W = 3.18 um; L = 2.00 um
* M5/M6: W = 1.57 um; L = 2.00 um
* M7/M8: W = 1.69 um; L = 2.00 um
* M9:    W = 38.21 um; L = 2.00 um
* M10:   W = 10.14 um; L = 2.00 um
* M11:   W = 6.37 um; L = 2.00 um
* M12:   W = 6.37 um; L = 2.00 um
* M13:   W = 1.69 um; L = 2.00 um
* M14:   W = 1.57 um; L = 2.00 um
* M15:   W = 1.57 um; L = 2.00 um
* IBIAS: 0.85 uA
* VIN MAX:   0.75 V
* VIN MIN:   -0.15 V
* VDSAT1:   0.10 V
* VIN:   0.30 V
* VOUT:  0.60 V
* Cf:    2.43 pF

*******************************

*** Supply voltage
.param vdd_val = 1.2

*** Load capacitance
.param Cl_val = 10p

*** Transistor dimensions

.param W1 = 3.18u
.param L1 = 2u
.param W2 = W1
.param L2 = L1

.param W3 = 3.18u
.param L3 = 2u
.param W4 = W3
.param L4 = L3

.param W5 = 1.57u
.param L5 = 2u
.param W6 = W5
.param L6 = 2u

.param W7 = 1.69u
.param L7 = 2u
.param W8 = W7
.param L8 = 2u

.param W9 = 38.21u
.param L9 = 2u
.param W10 = 10.14u
.param L10 = 2u
.param W11 = 6.37u
.param L11 = 2u
.param W12 = 6.37u
.param L12 = 2u
.param W13 = 1.69u
.param L13 = 2u
.param W14 = 1.57u
.param L14 = 2u
.param W15 = 1.57u
.param L15 = 2u

.param Cf_val = 2.43p

*** Bias point

.param VIN = 0.30
.param IBIAS = 0.85u

*** AC simulation parameters

.param V0 = 5m
.param fmin = 1
.param fmax = 1e9
.param ac_dec = 20

*******************************
*	Device under test
*******************************

***** Miller OTA

* Reminder
* xMN D G S B


* netlist : 
* M14 VBIAS2 VBIAS2 0 0 NMOS
* M13 VBIAS3 VBIAS2 0 0 NMOS
* M15 VBIAS1 VBIAS1 VBIAS2 VBIAS2 NMOS
* M7 N007 VBIAS2 0 0 NMOS
* M8 N006 VBIAS2 0 0 NMOS
* M6 N001 VBIAS1 N007 N007 NMOS
* M5 N002 VBIAS1 N006 N006 NMOS
* M10 N003 VBIAS2 0 0 NMOS
* C1 N003 N002 Cm
* C2 N003 0 CL
* M4 N001 N001 VDD VDD PMOS
* M3 N002 N001 VDD VDD PMOS
* M9 N003 N002 VDD VDD PMOS
* M2 N006 VIN+ N005 N005 PMOS
* M1 N007 VIN- N005 N005 PMOS
* M11 N005 VBIAS3 VDD VDD PMOS
* M12 VBIAS3 VBIAS3 VDD VDD PMOS
* I1 VDD VBIAS1 I

xM1 N007 INm N005 N005 pch_lvt_mac W=W1 L=L1
xM2 N006 INp N005 N005 pch_lvt_mac W=W2 L=L2

xM3 N002 N001 VDD VDD pch_lvt_mac W=W3 L=L3
xM4 N001 N001 VDD VDD pch_lvt_mac W=W4 L=L4
xM5 N002 VBIAS1 N006 N006 nch_lvt_mac W=W5 L=L5
xM6 N001 VBIAS1 N007 N007 nch_lvt_mac W=W6 L=L6

xM7 N007 VBIAS2 GND GND nch_lvt_mac W=W7 L=L7
xM8 N006 VBIAS2 GND GND nch_lvt_mac W=W8 L=L8

xM9 OUT N002 VDD VDD pch_lvt_mac W=W9 L=L9
xM10 OUT VBIAS2 GND GND nch_lvt_mac W=W10 L=L10

xM11 N005 VBIAS3 VDD VDD pch_lvt_mac W=W11 L=L11
xM12 VBIAS3 VBIAS3 VDD VDD pch_lvt_mac W=W12 L=L12

xM13 VBIAS3 VBIAS2 GND GND nch_lvt_mac W=W13 L=L13
xM14  VBIAS2 VBIAS2 GND GND nch_lvt_mac W=W14 L=L14
xM15 VBIAS1 VBIAS1 VBIAS2 VBIAS2 nch_lvt_mac W=W15 L=L15
Cf OUT N002 Cf_val

* Load capacitance
Cload OUT GND Cl_val
	
**********************************
*	Supply and stimuli
**********************************

*** Ideal current source	
IIbias VDD VBIAS1 DC IBIAS

*** Ground
* absolute voltage reference
.connect GND 0

*** Supply voltage
VVDD VDD GND DC vdd_val

*** Input Voltages Sources

***** DC & AC *****

VVINp INp GND DC VIN AC +V0
VVINm INm GND DC VIN AC -V0

**********************************
*	Simulations and Measurements
**********************************

***** DC *****

.OP

.extract DC label=IN V(INp)
.extract DC label=VOUT V(OUT)
.extract DC label=VSG12 -VGS(xM1.MAIN)
.extract DC label=VSD1 -VDS(xM1.MAIN)
.extract DC label=VSD2 -VDS(xM2.MAIN)
.extract DC label=VGS34 -VGS(xM3.MAIN)
.extract DC label=VDS3 -VDS(xM3.MAIN)
.extract DC label=VDS4 -VDS(xM4.MAIN)
.extract DC label=VGS5 VGS(xM5.MAIN)
.extract DC label=VDS5 VDS(xM5.MAIN)
.extract DC label=VSG6 VGS(xM6.MAIN)
.extract DC label=VSD6 VDS(xM6.MAIN)
.extract DC label=VSG7 VGS(xM7.MAIN)
.extract DC label=VSD7 VDS(xM7.MAIN)
.extract DC label=VSG8 VGS(xM8.MAIN)
.extract DC label=VSD8 VDS(xM8.MAIN)
.extract DC label=VSG9 -VGS(xM9.MAIN)
.extract DC label=VSD9 -VDS(xM9.MAIN)
.extract DC label=VGS10 VGS(xM10.MAIN)
.extract DC label=VDS10 VDS(xM10.MAIN)
.extract DC label=VSG11 -VGS(xM11.MAIN)
.extract DC label=VSD11 -VDS(xM11.MAIN)
.extract DC label=VSD12 -VDS(xM12.MAIN)
.extract DC label=VSG13 VGS(xM13.MAIN)
.extract DC label=VSD13 VDS(xM13.MAIN)
.extract DC label=VSG14 VGS(xM14.MAIN)
.extract DC label=VSD14 VDS(xM14.MAIN)
.extract DC label=VSG15 VGS(xM15.MAIN)
.extract DC label=VSD15 VDS(xM15.MAIN)

*** Currents
.extract DC label=ID1  I(xM1.MAIN.S)
.extract DC label=ID2  I(xM2.MAIN.S)
.extract DC label=ID3  I(xM3.MAIN.S)
.extract DC label=ID4  I(xM4.MAIN.S)
.extract DC label=ID5  I(xM5.MAIN.D)
.extract DC label=ID6  I(xM6.MAIN.D)
.extract DC label=ID7  I(xM7.MAIN.D)
.extract DC label=ID8  I(xM8.MAIN.D)
.extract DC label=ID9  I(xM9.MAIN.S)
.extract DC label=ID10 I(xM10.MAIN.D)
.extract DC label=ID11 I(xM11.MAIN.S)
.extract DC label=ID12 I(xM12.MAIN.S)
.extract DC label=ID13 I(xM13.MAIN.D)
.extract DC label=ID14 I(xM14.MAIN.D)
.extract DC label=ID15 I(xM15.MAIN.D)

* (gm/ID)'s 
.extract DC label=gm_over_ID1 'gm(xM1.MAIN)/ID1'
.extract DC label=gm_over_ID2 'gm(xM2.MAIN)/ID2'
.extract DC label=gm_over_ID3 'gm(xM3.MAIN)/ID3'
.extract DC label=gm_over_ID4 'gm(xM4.MAIN)/ID4'
.extract DC label=gm_over_ID6 'gm(xM6.MAIN)/ID6'
.extract DC label=gm_over_ID7 'gm(xM7.MAIN)/ID7'
.extract DC label=gm_over_ID8 'gm(xM8.MAIN)/ID8'
.extract DC label=gm_over_ID9 'gm(xM9.MAIN)/ID9'
.extract DC label=gm_over_ID10 'gm(xM10.MAIN)/ID10'
.extract DC label=gm_over_ID11 'gm(xM11.MAIN)/ID11'
.extract DC label=gm_over_ID12 'gm(xM12.MAIN)/ID12'
.extract DC label=gm_over_ID13 'gm(xM13.MAIN)/ID13'
.extract DC label=gm_over_ID14 'gm(xM14.MAIN)/ID14'
.extract DC label=gm_over_ID15 'gm(xM15.MAIN)/ID15'

* Power consumption
.extract DC label=Power 'V(VDD)*(-I(VVDD)-ID8)'

* Region of operation
.extract DC label=M1 opmode(xM1.MAIN)
.extract DC label=M2 opmode(xM2.MAIN)
.extract DC label=M3 opmode(xM3.MAIN)
.extract DC label=M4 opmode(xM4.MAIN)
.extract DC label=M5 opmode(xM5.MAIN)
.extract DC label=M6 opmode(xM6.MAIN)
.extract DC label=M7 opmode(xM7.MAIN)
.extract DC label=M8 opmode(xM8.MAIN)
.extract DC label=M9 opmode(xM9.MAIN)
.extract DC label=M10 opmode(xM10.MAIN)
.extract DC label=M11 opmode(xM11.MAIN)
.extract DC label=M12 opmode(xM12.MAIN)
.extract DC label=M13 opmode(xM13.MAIN)
.extract DC label=M14 opmode(xM14.MAIN)
.extract DC label=M15 opmode(xM15.MAIN)

***** AC *****


.AC dec ac_dec fmin fmax

*** Gain
.defwave Av = 'v(OUT)/(v(INp)-v(INm))'
.defwave Av1 = 'v(n1)/(v(INp)-v(INm))'
.defwave Av2 = 'v(OUT) / v(n1)'

.extract AC label=Av0 'max(wdb(Av))'
*** Transition Frequency
.extract AC label=fT 'xthres(wdb(Av),0)'
*** Phase Margin
.extract AC label=Phase_Margin '180 - yval(wp(Av),1) + xycond(wp(Av),wdb(Av)<0)'

*** Bode diagram (amplitude and phase)
.plot AC w(Av1) w(Av2)
.plot AC w(Av)